library IEEE;

use IEEE.std_logic_1164.all;

package divider_const is
	constant DIVIDEND_WIDTH : natural:= 8;
	constant DIVISOR_WIDTH : natural:= 4;
	
end package divider_const;

package body divider_const is
end package body divider_const;